LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY cw4 IS
PORT ( SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
HEX0 : OUT STD_LOGIC_VECTOR(0 TO 6);
HEX1 : OUT STD_LOGIC_VECTOR(0 TO 6);
HEX2 : OUT STD_LOGIC_VECTOR(0 TO 6);
HEX3 : OUT STD_LOGIC_VECTOR(0 TO 6);
HEX4 : OUT STD_LOGIC_VECTOR(0 TO 6);
HEX5 : OUT STD_LOGIC_VECTOR(0 TO 6);
HEX6 : OUT STD_LOGIC_VECTOR(0 TO 6);
HEX7 : OUT STD_LOGIC_VECTOR(0 TO 6));
END cw4;
ARCHITECTURE strukturalna OF cw4 IS
CONSTANT SPACJA: STD_LOGIC_VECTOR(2 DOWNTO 0):="000"; -- KOD SPACJI 
--DEKLARACJA KOMPONENTÓW
COMPONENT mux3bit_8to1 -- muliptekser
PORT ( S, U0, U1, U2, U3, U4, U5,U6,U7: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
--WEKTOR STERUJĄCY I 8 wektorów INFORMACYJNYCH
M0 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END COMPONENT;
COMPONENT char7seg -- transkoder
PORT (
 C : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
 Display : OUT STD_LOGIC_VECTOR(0 TO 6));
END COMPONENT;
SIGNAL M0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL M1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL M2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL M3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL M4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL M5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL M6 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL M7 : STD_LOGIC_VECTOR(2 DOWNTO 0);
 --do uzupełnienia
BEGIN
-- KONKRETYZACJA UŻYCIA KOMPONENTÓW
MUX0: mux3bit_8to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9),SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA,M0); 
MUX1: mux3bit_8to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9),SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA,M1);  
MUX2: mux3bit_8to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9),SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA,M2);  
MUX3: mux3bit_8to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9),SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA,M3);  
MUX4: mux3bit_8to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9),SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA,M4);  
MUX5: mux3bit_8to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9),SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA,M5);  
MUX6: mux3bit_8to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9),SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA,M6);   
MUX7: mux3bit_8to1 PORT MAP (SW(17 DOWNTO 15), SW(14 DOWNTO 12), SW(11 DOWNTO 9),SW(8 DOWNTO 6), SW(5 DOWNTO 3), SW(2 DOWNTO 0),SPACJA,SPACJA,SPACJA,M7);  

--do uzupełnienia
-- KONKRETYZACJE KOLEJNYCH MULTIPLEKSERÓW UKŁADU
H0: char7seg PORT MAP (M0, HEX0);
H1: char7seg PORT MAP (M1, HEX1);
H2: char7seg PORT MAP (M2, HEX2);
H3: char7seg PORT MAP (M3, HEX3);
H4: char7seg PORT MAP (M4, HEX4);
H5: char7seg PORT MAP (M5, HEX5);
H6: char7seg PORT MAP (M6, HEX6);
H7: char7seg PORT MAP (M7, HEX7);

--do uzupełnienia
-- KONKRETYZACJE KOLEJNYCH TRANSKODERÓW
END strukturalna;
-- implementacja multipleksera 8 do 1 (wektor 3 bitowy)
LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY mux3bit_8to1 IS 
PORT ( S, U0, U1, U2, U3, U4, U5,U6,U7: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
M0 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END mux3bit_8to1;
ARCHITECTURE strukturalna OF mux3bit_8to1 IS
Begin 
With S select 
M0 	<=	U0 when "000",
		U1 when "001",
		U2 when "010",
		U3 when "011",
		U4 when "100",
		U5 when "101",
		U6 when "110",
		U7 when "111";
-- do uzupełnienia
END strukturalna;
-- IMPLEMENTACJA TRANSKODERA
LIBRARY ieee;
USE ieee.std_logic_1164.all;
ENTITY char7seg IS
PORT ( C : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
Display : OUT STD_LOGIC_VECTOR(0 TO 6));
END char7seg;
ARCHITECTURE strukturalna OF char7seg IS
Begin
With C select Display <=
"0000000" when "000", --spacja
"0000110" when "001", -- I
"0111100" when "010", -- J
"0001110" when "011", -- L
"1111110" when "100", -- O
"0000000" when others;
-- douzupełnienia
END strukturalna;